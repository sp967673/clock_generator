//#
//#
//#

//# The CLK_UVC_FREQ_MHZ is used to define the reqiured clock frequency used in TB. Default value is 100 (100MHz)
`define CLK_UVC_FREQ_MHZ   100

//# The CLK_UVC_DUTY_CYCLE can use to select the frequency-specified duty cycle. Default value is 0.5 (50%)
`define CLK_UVC_DUTY_CYCLE 0.5

//# 
`define CLK_UVC_JITTER_MAX 5
`define CLK_UVC_JITTER_MIN 1
